// Company: uth university school of engineers
// Engineer: Dimkou Eleni
// 			 Karagiannis Marios
// 			 Lianidis Theodoros 
`timescale 1ns/1ps
`define clock_period  10

/*in_pc*/


module finaltb;

    reg clk;
    reg  [31:0] x1, y1, z1, x2, y2, z2, w1, w2;
    wire [31:0] length;
    wire [31:0] innerproduct;
    reg [3:0] func;
    wire [7:0] overflow;

    calculator calc (clk, x1, y1, z1, w1, x2, y2, z2, w2, length, innerproduct, func, overflow);

    initial   $dumpfile("final.vcd");
    initial   $dumpvars(0, finaltb);

    always #(`clock_period / 2) clk = ~clk;

    initial begin


		x1 = 0; y1 = 0; z1 = 0; w1 = 0;
        x2 = 0; y2 = 0; z2 = 0; w2 = 0;
		clk = 0;
        func = 4'b0000; //idle calc

        
        //$readmemb("program.txt", data, 0, 95);
		#200

        x1 = 32'b0000_0000_0000_0001_0000_0000_0000_0000; // 1
        y1 = 32'b0000_0000_0000_0010_0000_0000_0000_0000; // 2
        z1 = 32'b0000_0000_0000_0001_0000_0000_0000_0000; // 1
        w1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;// 0
        x2 = 32'b0000_0000_0000_0000_1000_0000_0000_0000; // 1/2
        y2 = 32'b0000_0000_0000_0101_0000_0000_0000_0000; // 5
        z2 = 32'b0000_0000_0000_0001_0000_0000_0000_0000; // 1
        w2 = 32'b0000_0000_0000_0001_1000_0000_0000_0000; // 1.5

        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

        x1 = 32'b0000_0000_0000_0000_0000_0000_1000_0000; // 0.003890
        y1 = 32'b1000_0000_0000_1100_0000_0000_0000_0000; // 0.98090
        z1 = 32'b0000_0000_0000_0000_1000_0000_0000_0000;// 0.5
        w1 = 32'b1000_0000_0000_0000_0100_0000_0000_0000; // -0.25
        x2 = 32'b0000_0000_0000_0001_1100_0000_0000_0000; // 1.75
        y2 = 32'b1000_0000_0000_0001_0000_0000_0000_0000; // -1
        z2 = 32'b1000_0000_0000_0001_0000_0000_0000_0000; // -1
        w2 = 32'b0000_0000_0000_0000_1000_0000_0000_0000; // 0.75

        
        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

            x1 = 32'b0000_0000_0000_0001_0000_0000_0000_0000; // 1
            y1 = 32'b0000_0000_0000_0001_0000_0000_0000_0000;
            z1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
            w1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
            x2 = 32'b0000_0000_0000_0001_1000_0000_0000_0000; // 1.5
            y2 = 32'b0000_0000_0000_0001_1000_0000_0000_0000;
            z2 = 32'b0000_0000_0000_0000_1000_0000_0000_0000; // 0.5
            w2 = 32'b0000_0000_0000_0010_0000_0000_0000_0000; // 2

            
        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

            x1 = 32'b1000_0000_0000_0001_0000_0000_0000_0000; // -1
            y1 = 32'b1000_0000_0000_0001_0000_0000_0000_0000;
            z1 = 32'b1000_0000_0000_0000_0110_0000_0000_0000; // 0.375
            w1 = 32'b1000_0000_0000_0000_0000_0000_0000_0000; // 0
            x2 = 32'b1000_0000_0000_0001_1000_0000_0000_0000; // -1.5
            y2 = 32'b1000_0000_0000_0001_1000_0000_0000_0000;
            z2 = 32'b1000_0000_0000_0000_1000_0000_0000_0000; // -0.5
            w2 = 32'b1000_0000_0000_0000_1000_0000_0000_0000;

            
        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

            x1 = 32'b0000_0000_0000_0001_0000_0000_0000_0000; // 1
            y1 = 32'b0000_0000_0000_0000_1000_0000_0000_0000;// 0.5
            z1 = 32'b1000_0000_0000_0001_0000_0000_0000_0000; // -1
            w1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
            x2 = 32'b0000_0000_0000_0001_0000_0000_0000_0000; // 1
            y2 = 32'b0000_0000_0000_0001_0000_0000_0000_0000; // 1
            z2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
            w2 = 32'b0000_0000_0000_0010_0000_0000_0000_0000; // 2

           
        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

            x1 = 32'b0000_0000_0001_0000_0000_0000_0000_0000; // 16
            y1 = 32'b0000_0000_0000_1100_0000_0000_0000_0000; // 12
            z1 = 32'b0000_0000_0000_0100_0000_0000_0000_0000; // 4
            w1 = 32'b1000_0000_0000_0001_0000_0000_0000_0000;// -1
            x2 = 32'b0000_0000_0000_0001_0000_0000_0000_0000; // 1
            y2 = 32'b1000_0000_0000_0001_0000_0000_0000_0000; // -1
            z2 = 32'b1000_0000_0000_0001_0000_0000_0000_0000; // -1
            w2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
            
            
        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

            x1 = 32'b0000_0000_0001_0000_1001_0000_0000_0000;// 16.5625
            y1 = 32'b0000_0000_0000_1100_0101_0100_0100_0000; // 12.3291
            z1 = 32'b0000_0000_0000_0100_1110_0100_1000_0000; // 4.89257
            w1 = 32'b1000_0000_0000_0001_1000_0000_0000_0000; // -1.5
            x2 = 32'b0000_0000_0000_0001_1111_1100_0000_0000; // 1.98090
            y2 = 32'b1000_0000_0000_0011_0000_0000_0000_0000; // -3
            z2 = 32'b1000_0000_0000_1001_0000_0000_0000_0000; // -9
            w2 = 32'b0000_0000_0000_0000_0000_0000_1111_1111; // 0.003890

            
        #1000 func = 4'b0000; //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

            x1 = 32'b0000_0000_0001_0100_0000_0000_0000_0000; // 20
            y1 = 32'b0000_0000_0000_1000_0000_0000_0000_0000; // 8
            z1 = 32'b1000_0000_0000_0100_0000_0000_0000_0000; // -4
            w1 = 32'b0000_0000_0001_1001_0000_0000_0000_0000; // 25
            x2 = 32'b1000_0000_0000_1001_0000_0000_0000_0000; // -9
            y2 = 32'b1000_0000_0000_0001_1000_0000_0000_0000; // -1.5
            z2 = 32'b1000_0000_0000_1010_0000_0000_0000_0000; // -10
            w2 = 32'b0000_0000_0000_0000_0000_1010_0000_0000; // 0.4 = 0.0390625

            
        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

            x1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
            y1 = 32'b0110_0000_0001_0010_0000_0000_0000_0000; // -32768  // FAULT sto mul gia length
            z1 = 32'b0000_0000_0000_0000_0011_0000_0011_0000; // 0.249969
            w1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;// 0
            x2 = 32'b0000_0000_0000_0000_0000_0000_0000_0010; // 0.000030517
            y2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
            z2 = 32'b0000_0000_0000_0100_0100_0000_0000_0000; // 4.25
            w2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0

           
        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

        x1 = 32'b0000_0000_0110_0100_0000_0000_0000_0000; // 100
        y1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
        z1 = 32'b0000_0000_1001_0110_0000_0000_0000_0000;// 150
        w1 = 32'b0000_0000_0001_0000_0000_0000_0000_0000; // 16
        x2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;// 0
        y2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
        z2 = 32'b0000_0000_0000_0001_0000_0000_0000_0000; // 1
        w2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0

            
        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

        x1 = 32'b1000_0000_1011_0100_1111_1100_0000_0000; // -180.984375
        y1 = 32'b0000_0000_0000_0010_0000_0000_0000_0000;// 2
        z1 = 32'b1000_0000_0001_0000_0000_0000_0000_0000; // -16
        w1 = 32'b0000_0000_0001_0000_0000_0000_0000_0000; // 0
        x2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
        y2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
        z2 = 32'b1000_0000_0000_0001_0010_0000_0000_0000; // -1.125
        w2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0

            
        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b1111; //4d inner product
        #1000 func = 4'b0000;
        #1000

        x1 = 32'b0000_0000_1000_0001_0000_0000_0000_0000; // 129  FAULT sto sum
        y1 = 32'b0000_0000_1000_0000_0000_0000_0000_0000;// 128
        z1 = 32'b0000_0000_0000_0010_0000_0000_0000_0000; // 2
        w1 = 32'b0000_0000_0000_0000_0001_0000_0000_0000; // 0.0625 1/16
        x2 = 32'b0000_0000_0000_0000_0000_0010_0000_0000; // 1/128
        y2 = 32'b0000_0000_0000_0010_0000_0000_0000_0000; // 2
        z2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000; // 0
        w2 = 32'b0000_0000_0001_0000_0000_0000_0000_0000;// 16

        #1000 func = 4'b1000;  //2d length
        #1000 func = 4'b1010; //3d length
        #1000 func = 4'b1011; //4d length
        #1000 func = 4'b1100; //2d inner product
        #1000 func = 4'b1110; //3d inner product
        #1000 func = 4'b0000; //4d inner product
        #1000 func = 4'b0000;
        #1000
         

		#25000 $finish;
		end
endmodule
